module teste;
integer A, B, C;
initial begin
A = 0;
B = 4;
C = 5;
$display("Here's your numbers -> %d, %d, %d", A, B, C);
end
endmodule