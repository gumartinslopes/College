module HelloWorld;
initial begin
    $display("Hello World I am on verilog");
end
endmodule